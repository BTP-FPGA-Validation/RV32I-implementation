e
 // Control Unit
module Control_Unit(instruction, Branch, MemRead, MemtoReg, ALUOp, MemWrite, ALUSrc, RegWrite);
 input [6:0] instruction;
 output reg Branch, MemRead, MemtoReg, MemWrite, ALUSrc, RegWrite;
 output reg [1:0] ALUOp;
always @(*) begin
  case (instruction)
    7'b0110011: begin // R-type
      ALUSrc   <= 0;
      MemtoReg <= 0;
      RegWrite <= 1;
      MemRead  <= 0;
      MemWrite <= 0;
      Branch   <= 0;
      ALUOp    <= 2'b10;
    end

    7'b0010011: begin // I-type (ADDI, ORI, etc.)
      ALUSrc   <= 1;
      MemtoReg <= 0;
      RegWrite <= 1;   // enable write
      MemRead  <= 0;
      MemWrite <= 0;
      Branch   <= 0;
      ALUOp    <= 2'b10;
    end

    7'b0000011: begin // Load
      ALUSrc   <= 1;
      MemtoReg <= 1;
      RegWrite <= 1;
      MemRead  <= 1;
      MemWrite <= 0;
      Branch   <= 0;
      ALUOp    <= 2'b00;
    end

    7'b0100011: begin // Store
      ALUSrc   <= 1;
      MemtoReg <= 0;
      RegWrite <= 0;
      MemRead  <= 0;
      MemWrite <= 1;
      Branch   <= 0;
      ALUOp    <= 2'b00;
    end

    7'b1100011: begin // Branch
      ALUSrc   <= 0;
      MemtoReg <= 0;
      RegWrite <= 0;
      MemRead  <= 0;
      MemWrite <= 0;
      Branch   <= 1;
      ALUOp    <= 2'b01;
    end

    default: begin
      ALUSrc   <= 0;
      MemtoReg <= 0;
      RegWrite <= 0;
      MemRead  <= 0;
      MemWrite <= 0;
      Branch   <= 0;
      ALUOp    <= 2'b00;
    end
  endcase
end


endmodule

